module InstructionMemory (
    input [4:0] Address,    // 5-bit address input to select one of 32 instructions
    output reg [31:0] Instruction  // 32-bit instruction output
);

    // Define a distributed RAM with 32 32-bit instructions
    reg [31:0] memory [31:0];
        // memory[0] = 32'b000000000011_00001_000_00010_0010011; // addi r2, r1, 3
        // memory[1] = 32'b000000000001_00001_000_00001_0010011; // addi r2, r1, 1
        // memory[2] = 32'b11111110001000001001111011100011; // bne r1, r2, -8
    // Initialize the instructions
    initial begin
        memory[0]  = 32'bx; // addi r0, r1, 3  (r2 = rb1 + 3)
        memory[1]  = 32'b00000000000100000000000110010011; // addi r3, r2, 1  (r3 = r2 + 1)
        memory[2]  = 32'b00000000001100000010000110100011; // sw r3, 3(r0)    (memory[r0 + 3] = r3)
        memory[3]  = 32'b00000000001100000010001000000011; // lw r4, 3(r0)    (r4 = memory[r0 + 3])
        memory[4]  = 32'b000000000000_00100_000_00001_1100011; // beq r4, r0, 4   (if r4 == r0, PC += 4)
        memory[5]  = 32'b00000000001100000010000110100011; // addi r1, r1, -1 (r1 = r1 - 1)
        memory[6]  = 32'b00000000001100000010001000000011; // addi r2, r2, 1  (r2 = r2 + 1)
        memory[7]  = 32'b111111111111_00001_000_00001_1100011; // bne r1, r0, -8  (if r1 != r0, PC -= 8)
        memory[8]   =32'b000000000011_00001_000_00010_0010011; // addi r2, r1, 3
        memory[9]   =32'b000000000001_00001_000_00001_0010011; // addi r2, r1, 1
        memory[10]   =32'b11111110001000001001111011100011; // bne r1, r2, -8
                // // // R        mtructions (addemory[16] = ; // add r3, r1, r2
        // memory[9]  =  32'b000000000011_00001_000_00010_0010011; // addi r2, r1, 3
        // memory[10] =  32'b000000000001_00001_000_00001_0010011; // addi r2, r1, 1
        // memory[19] =  32'b11111110001000001001111011100011; // bne r1, r2, -8
        // memory[20] = 32'b0100000_00111_01000_000_01001_0110011; // add r11, r9, r10
        // memory[21] = 32'b0000000_01001_01010_000_01011_0110011; // sub r13, r11, r12
        // memory[22] = 32'b0100000_01011_01100_000_01101_0110011; // add r15, r13, r14
        // memory[23] = 32'b0000000_01101_01110_000_01111_0110011; // sub r17, r15, r16
        // memory[24] = 32'b0100000_01111_10000_000_10001_0110011; // add r19, r17, r18
        // memory[25] = 32'b0000000_10001_10010_000_10011_0110011; // sub r21, r19, r20
        // memory[26] = 32'b0100000_10011_10100_000_10101_0110011; // add r23, r21, r22
        // memory[27] = 32'b0000000_10101_10110_000_10111_0110011; // sub r25, r23, r24
        // memory[28] = 32'b0100000_10111_11000_000_11001_0110011; // add r27, r25, r26
        // memory[29] = 32'b0000000_11001_11010_000_11011_0110011; // sub r29, r27, r28
        // memory[30] = 32'b0100000_11011_11100_000_11101_0110011; // add r31, r29, r30
        // memory[31] = 32'b0000000_11101_11110_000_11111_0110011; // sub r1, r31, r0
    end

    // Read instruction based on address
    always @(*) begin
        Instruction = memory[Address];
    end

endmodule
